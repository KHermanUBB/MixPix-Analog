** sch_path: /home/icarosix/asic/MixPix/MixPix-Analog/xchem/OTA3_lvt.sch
**.subckt OTA3_lvt
C1 Vout GND 20f m=1
V2 VDD GND 1.8
V1 Vin_p net1 dc 0 ac 0.1m sin(0 100u 50)
V3 Vin_n net2 dc 0 ac 0 sin(0 -100u 50)
V4 net1 GND 0.9
V5 net2 GND 0.9
XM1 Vas Vin_n Vsrc GND sky130_fd_pr__nfet_01v8_lvt L=1 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vmid Vin_p Vsrc GND sky130_fd_pr__nfet_01v8_lvt L=1 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 Vas Vas VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 Vmid Vas VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 Vout Vmid VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=5.1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 Vout Vcs GND GND sky130_fd_pr__nfet_01v8_lvt L=1 W=2.90 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 Vsrc Vcs GND GND sky130_fd_pr__nfet_01v8_lvt L=0.5 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 Vcs Vcs GND GND sky130_fd_pr__nfet_01v8_lvt L=0.5 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 Vcs net3 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
C2 Vout Vmid 300f m=1
XM10 net3 net3 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.8 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM11 net3 net4 GND GND sky130_fd_pr__nfet_01v8_lvt L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM12 net4 net4 GND GND sky130_fd_pr__nfet_01v8_lvt L=0.5 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
I0 GND net4 120u
**** begin user architecture code


.control
run
save all
*tran 10u 100m
*plot Vout
ac dec 101 1 1g
plot db(1*V(Vout)/(V(Vin_p) - V(Vin_n))), 180/PI*phase(V(Vout))


let id1  = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[id]
let id2  = @m.xm2.msky130_fd_pr__nfet_01v8_lvt[id]
let id3  = @m.xm3.msky130_fd_pr__pfet_01v8_lvt[id]
let id4  = @m.xm4.msky130_fd_pr__pfet_01v8_lvt[id]
let id5  = @m.xm5.msky130_fd_pr__pfet_01v8_lvt[id]
let id6  = @m.xm6.msky130_fd_pr__nfet_01v8_lvt[id]
let id7  = @m.xm7.msky130_fd_pr__nfet_01v8_lvt[id]
let id8  = @m.xm8.msky130_fd_pr__nfet_01v8_lvt[id]

let gm1  = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
let gm2  = @m.xm2.msky130_fd_pr__nfet_01v8_lvt[gm]
let gm3  = @m.xm3.msky130_fd_pr__pfet_01v8_lvt[gm]
let gm4  = @m.xm4.msky130_fd_pr__pfet_01v8_lvt[gm]
let gm5  = @m.xm5.msky130_fd_pr__pfet_01v8_lvt[gm]
let gm6  = @m.xm6.msky130_fd_pr__nfet_01v8_lvt[gm]
let gm7  = @m.xm7.msky130_fd_pr__nfet_01v8_lvt[gm]
let gm8  = @m.xm8.msky130_fd_pr__nfet_01v8_lvt[gm]

let gds1  = @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gds]
let gds2  = @m.xm2.msky130_fd_pr__nfet_01v8_lvt[gds]
let gds3  = @m.xm3.msky130_fd_pr__pfet_01v8_lvt[gds]
let gds4  = @m.xm4.msky130_fd_pr__pfet_01v8_lvt[gds]
let gds5  = @m.xm5.msky130_fd_pr__pfet_01v8_lvt[gds]
let gds6  = @m.xm6.msky130_fd_pr__nfet_01v8_lvt[gds]

let Av1  = gm2/(gds2+gds4)
let Av2  = gm5/(gds5 + gds6)
let Av = Av1*Av2

let Cl = 20e-15
let Cn5 = @m.xm5.msky130_fd_pr__pfet_01v8_lvt[cgs]
let GBW = gm1/(6.28*(Cl + Cn5))

print gm1/id1
print gm2/id2
print gm3/id3
print gm4/id4
print gm5/id5
print gm6/id6
print gm7/id7
print gm8/id8

print Av1
print Av2
print Av
print GBW

.endc



** opencircuitdesign pdks install
.lib /home/icarosix/asic/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends
.GLOBAL GND
.end
