magic
tech sky130A
magscale 1 2
timestamp 1663448264
<< nwell >>
rect -683 -312 683 312
<< pmoslvt >>
rect -487 -92 -287 164
rect -229 -92 -29 164
rect 29 -92 229 164
rect 287 -92 487 164
<< pdiff >>
rect -545 152 -487 164
rect -545 -80 -533 152
rect -499 -80 -487 152
rect -545 -92 -487 -80
rect -287 152 -229 164
rect -287 -80 -275 152
rect -241 -80 -229 152
rect -287 -92 -229 -80
rect -29 152 29 164
rect -29 -80 -17 152
rect 17 -80 29 152
rect -29 -92 29 -80
rect 229 152 287 164
rect 229 -80 241 152
rect 275 -80 287 152
rect 229 -92 287 -80
rect 487 152 545 164
rect 487 -80 499 152
rect 533 -80 545 152
rect 487 -92 545 -80
<< pdiffc >>
rect -533 -80 -499 152
rect -275 -80 -241 152
rect -17 -80 17 152
rect 241 -80 275 152
rect 499 -80 533 152
<< nsubdiff >>
rect -647 242 -551 276
rect 551 242 647 276
rect -647 179 -613 242
rect 613 179 647 242
rect -647 -242 -613 -179
rect 613 -242 647 -179
rect -647 -276 -551 -242
rect 551 -276 647 -242
<< nsubdiffcont >>
rect -551 242 551 276
rect -647 -179 -613 179
rect 613 -179 647 179
rect -551 -276 551 -242
<< poly >>
rect -487 164 -287 190
rect -229 164 -29 190
rect 29 164 229 190
rect 287 164 487 190
rect -487 -139 -287 -92
rect -487 -173 -471 -139
rect -303 -173 -287 -139
rect -487 -189 -287 -173
rect -229 -139 -29 -92
rect -229 -173 -213 -139
rect -45 -173 -29 -139
rect -229 -189 -29 -173
rect 29 -139 229 -92
rect 29 -173 45 -139
rect 213 -173 229 -139
rect 29 -189 229 -173
rect 287 -139 487 -92
rect 287 -173 303 -139
rect 471 -173 487 -139
rect 287 -189 487 -173
<< polycont >>
rect -471 -173 -303 -139
rect -213 -173 -45 -139
rect 45 -173 213 -139
rect 303 -173 471 -139
<< locali >>
rect -647 242 -551 276
rect 551 242 647 276
rect -647 179 -613 242
rect 613 179 647 242
rect -533 152 -499 168
rect -533 -96 -499 -80
rect -275 152 -241 168
rect -275 -96 -241 -80
rect -17 152 17 168
rect -17 -96 17 -80
rect 241 152 275 168
rect 241 -96 275 -80
rect 499 152 533 168
rect 499 -96 533 -80
rect -487 -173 -471 -139
rect -303 -173 -287 -139
rect -229 -173 -213 -139
rect -45 -173 -29 -139
rect 29 -173 45 -139
rect 213 -173 229 -139
rect 287 -173 303 -139
rect 471 -173 487 -139
rect -647 -242 -613 -179
rect 613 -242 647 -179
rect -647 -276 -551 -242
rect 551 -276 647 -242
<< viali >>
rect -533 -80 -499 152
rect -275 -80 -241 152
rect -17 -80 17 152
rect 241 -80 275 152
rect 499 -80 533 152
rect -471 -173 -303 -139
rect -213 -173 -45 -139
rect 45 -173 213 -139
rect 303 -173 471 -139
<< metal1 >>
rect -539 152 -493 164
rect -539 -80 -533 152
rect -499 -80 -493 152
rect -539 -92 -493 -80
rect -281 152 -235 164
rect -281 -80 -275 152
rect -241 -80 -235 152
rect -281 -92 -235 -80
rect -23 152 23 164
rect -23 -80 -17 152
rect 17 -80 23 152
rect -23 -92 23 -80
rect 235 152 281 164
rect 235 -80 241 152
rect 275 -80 281 152
rect 235 -92 281 -80
rect 493 152 539 164
rect 493 -80 499 152
rect 533 -80 539 152
rect 493 -92 539 -80
rect -483 -139 -291 -133
rect -483 -173 -471 -139
rect -303 -173 -291 -139
rect -483 -179 -291 -173
rect -225 -139 -33 -133
rect -225 -173 -213 -139
rect -45 -173 -33 -139
rect -225 -179 -33 -173
rect 33 -139 225 -133
rect 33 -173 45 -139
rect 213 -173 225 -139
rect 33 -179 225 -173
rect 291 -139 483 -133
rect 291 -173 303 -139
rect 471 -173 483 -139
rect 291 -179 483 -173
<< properties >>
string FIXED_BBOX -630 -259 630 259
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.28 l 1.0 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
