magic
tech sky130A
magscale 1 2
timestamp 1663456995
<< nwell >>
rect -4020 2850 -300 3660
rect -4020 2760 -275 2850
rect -4000 2088 -2725 2275
rect -2250 2000 -1900 2760
rect -1350 2508 -275 2760
<< locali >>
rect -3798 3030 -3672 3234
rect -3156 3030 -2754 3234
rect -2898 3024 -2754 3030
rect -1296 2958 -1248 3072
rect -780 2958 -732 3060
rect -4062 2784 -342 2958
rect -2350 2775 -1900 2784
rect -3798 2676 -2376 2718
rect -1884 2676 -474 2718
rect -2350 2025 -1900 2075
rect -3348 1776 -804 1824
rect -3708 1362 -3570 1638
rect -690 1584 -540 1680
rect -696 1578 -540 1584
rect -696 1302 -420 1578
rect -4068 1152 -3564 1212
rect -3396 1152 -3360 1248
rect -2880 1152 -2844 1248
rect -2364 1152 -2328 1248
rect -1848 1152 -1812 1260
rect -1332 1152 -1296 1260
rect -804 1212 -768 1260
rect -696 1212 -540 1302
rect -804 1152 -144 1212
rect -4068 1092 -144 1152
rect -4068 1086 -3936 1092
<< metal1 >>
rect -1482 3414 -546 3450
rect -3642 3312 -2550 3318
rect -1482 3312 -1446 3414
rect -3642 3276 -1446 3312
rect -3456 2988 -3384 3228
rect -4062 2928 -3384 2988
rect -4062 2922 -3390 2928
rect -4062 2916 -3396 2922
rect -4062 2910 -3996 2916
rect -2532 2856 -2472 3240
rect -1032 2988 -996 3072
rect -516 2988 -480 3072
rect -1032 2940 -48 2988
rect -132 2916 -48 2940
rect -3552 2814 -720 2856
rect -3558 2778 -720 2814
rect -3912 2088 -3840 2628
rect -3558 2616 -3516 2778
rect -2958 2616 -2916 2778
rect -2580 2736 -2400 2748
rect -2580 2676 -2568 2736
rect -2412 2676 -2400 2736
rect -2580 2664 -2400 2676
rect -2364 2616 -2322 2778
rect -1956 2604 -1914 2778
rect -1884 2676 -1872 2748
rect -1692 2676 -1680 2748
rect -1356 2610 -1314 2778
rect -762 2610 -720 2778
rect -3252 2088 -3216 2160
rect -2652 2088 -2616 2184
rect -1656 2100 -1614 2184
rect -1062 2100 -1020 2184
rect -462 2100 -420 2190
rect -3912 2052 -2616 2088
rect -3912 1728 -3840 2052
rect -1668 2028 -228 2100
rect -3774 1884 -339 1926
rect -3774 1728 -3732 1884
rect -1020 1818 -804 1824
rect -1020 1764 -990 1818
rect -828 1764 -804 1818
rect -1020 1758 -804 1764
rect -3912 1680 -3732 1728
rect -3912 1572 -3840 1680
rect -381 1623 -339 1884
rect -288 1824 -228 2028
rect -306 1818 -162 1824
rect -306 1764 -294 1818
rect -306 1758 -162 1764
rect -3912 1344 -3852 1572
rect -288 1284 -228 1758
rect -3138 1176 -3096 1260
rect -2622 1176 -2580 1260
rect -2106 1176 -2064 1260
rect -1590 1176 -1548 1260
rect -1074 1176 -1032 1260
rect -132 1176 -72 2916
rect -3138 1092 -72 1176
<< via1 >>
rect -2568 2676 -2412 2736
rect -1872 2676 -1692 2748
rect -990 1764 -828 1818
rect -294 1764 -162 1818
<< metal2 >>
rect -4068 3480 -2256 3552
rect -4068 3372 -2364 3444
rect -2436 2748 -2364 3372
rect -2580 2736 -2364 2748
rect -2580 2676 -2568 2736
rect -2412 2676 -2364 2736
rect -2328 2748 -2256 3480
rect -1896 2748 -1668 2760
rect -2328 2676 -1872 2748
rect -1692 2676 -1668 2748
rect -2580 2664 -2400 2676
rect -1896 2664 -1668 2676
rect -1068 1824 -780 1848
rect -1068 1752 -1044 1824
rect -804 1818 -150 1824
rect -804 1764 -294 1818
rect -162 1764 -150 1818
rect -804 1758 -150 1764
rect -804 1752 -780 1758
rect -1068 1728 -780 1752
<< via2 >>
rect -1044 1818 -804 1824
rect -1044 1764 -990 1818
rect -990 1764 -828 1818
rect -828 1764 -804 1818
rect -1044 1752 -804 1764
<< metal3 >>
rect -1572 2988 -1440 3072
rect -1500 1824 -1440 2988
rect -1068 1824 -780 1848
rect -1500 1764 -1044 1824
rect -1068 1752 -1044 1764
rect -804 1752 -780 1824
rect -1068 1728 -780 1752
use sky130_fd_pr__pfet_01v8_lvt_UXWVYC  XM2
timestamp 1663451206
transform 1 0 -3088 0 1 2424
box -912 -424 912 424
use sky130_fd_pr__nfet_01v8_lvt_9MXGXM  XM3
timestamp 1663453301
transform 1 0 -353 0 1 1470
box -246 -329 246 329
use sky130_fd_pr__nfet_01v8_lvt_PVELEM  XM4
timestamp 1663448021
transform 1 0 -3774 0 1 1500
box -246 -360 246 360
use sky130_fd_pr__pfet_01v8_lvt_P7LFVU  XM5
timestamp 1663453301
transform 1 0 -886 0 1 3235
box -554 -355 554 355
use sky130_fd_pr__nfet_01v8_lvt_E8GDTS  XM6
timestamp 1663448045
transform 1 0 -2083 0 1 1509
box -1457 -429 1457 429
use sky130_fd_pr__pfet_01v8_lvt_SPR9VP  XM7
timestamp 1663449709
transform 1 0 -2644 0 1 3164
box -296 -284 296 284
use sky130_fd_pr__pfet_01v8_lvt_7PHJSE  XM8
timestamp 1663449709
transform 1 0 -3415 0 1 3164
box -425 -284 425 284
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_0
timestamp 1663456995
transform 1 0 -1846 0 1 3228
box -350 -300 349 300
use sky130_fd_pr__pfet_01v8_lvt_UXWVYC  sky130_fd_pr__pfet_01v8_lvt_UXWVYC_0
timestamp 1663451206
transform 1 0 -1188 0 1 2424
box -912 -424 912 424
<< labels >>
flabel metal2 -4068 3408 -4068 3408 0 FreeSans 80 0 0 0 IN_M
port 1 nsew
flabel metal2 -4068 3516 -4068 3516 0 FreeSans 80 0 0 0 IN_P
port 2 nsew
flabel metal1 -4056 2976 -4056 2976 0 FreeSans 80 0 0 0 Ib
port 3 nsew
flabel locali -4056 2868 -4056 2868 0 FreeSans 80 0 0 0 VCC
port 5 nsew
flabel locali -4056 1152 -4056 1152 0 FreeSans 80 0 0 0 GND
port 6 nsew
flabel metal1 -60 2952 -60 2952 0 FreeSans 80 0 0 0 Out
port 7 nsew
<< end >>
