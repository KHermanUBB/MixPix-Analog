magic
tech sky130A
magscale 1 2
timestamp 1663450919
<< nwell >>
rect -912 -424 912 424
<< pmoslvt >>
rect -716 -276 -476 204
rect -418 -276 -178 204
rect -120 -276 120 204
rect 178 -276 418 204
rect 476 -276 716 204
<< pdiff >>
rect -774 192 -716 204
rect -774 -264 -762 192
rect -728 -264 -716 192
rect -774 -276 -716 -264
rect -476 192 -418 204
rect -476 -264 -464 192
rect -430 -264 -418 192
rect -476 -276 -418 -264
rect -178 192 -120 204
rect -178 -264 -166 192
rect -132 -264 -120 192
rect -178 -276 -120 -264
rect 120 192 178 204
rect 120 -264 132 192
rect 166 -264 178 192
rect 120 -276 178 -264
rect 418 192 476 204
rect 418 -264 430 192
rect 464 -264 476 192
rect 418 -276 476 -264
rect 716 192 774 204
rect 716 -264 728 192
rect 762 -264 774 192
rect 716 -276 774 -264
<< pdiffc >>
rect -762 -264 -728 192
rect -464 -264 -430 192
rect -166 -264 -132 192
rect 132 -264 166 192
rect 430 -264 464 192
rect 728 -264 762 192
<< nsubdiff >>
rect -876 354 -780 388
rect 780 354 876 388
rect -876 291 -842 354
rect 842 291 876 354
rect -876 -354 -842 -291
rect 842 -354 876 -291
rect -876 -388 -780 -354
rect 780 -388 876 -354
<< nsubdiffcont >>
rect -780 354 780 388
rect -876 -291 -842 291
rect 842 -291 876 291
rect -780 -388 780 -354
<< poly >>
rect -716 285 -476 301
rect -716 251 -700 285
rect -492 251 -476 285
rect -716 204 -476 251
rect -418 285 -178 301
rect -418 251 -402 285
rect -194 251 -178 285
rect -418 204 -178 251
rect -120 285 120 301
rect -120 251 -104 285
rect 104 251 120 285
rect -120 204 120 251
rect 178 285 418 301
rect 178 251 194 285
rect 402 251 418 285
rect 178 204 418 251
rect 476 285 716 301
rect 476 251 492 285
rect 700 251 716 285
rect 476 204 716 251
rect -716 -302 -476 -276
rect -418 -302 -178 -276
rect -120 -302 120 -276
rect 178 -302 418 -276
rect 476 -302 716 -276
<< polycont >>
rect -700 251 -492 285
rect -402 251 -194 285
rect -104 251 104 285
rect 194 251 402 285
rect 492 251 700 285
<< locali >>
rect -876 354 -780 388
rect 780 354 876 388
rect -876 291 -842 354
rect 842 291 876 354
rect -716 251 -700 285
rect -492 251 -476 285
rect -418 251 -402 285
rect -194 251 -178 285
rect -120 251 -104 285
rect 104 251 120 285
rect 178 251 194 285
rect 402 251 418 285
rect 476 251 492 285
rect 700 251 716 285
rect -762 192 -728 208
rect -762 -280 -728 -264
rect -464 192 -430 208
rect -464 -280 -430 -264
rect -166 192 -132 208
rect -166 -280 -132 -264
rect 132 192 166 208
rect 132 -280 166 -264
rect 430 192 464 208
rect 430 -280 464 -264
rect 728 192 762 208
rect 728 -280 762 -264
rect -876 -354 -842 -291
rect 842 -354 876 -291
rect -876 -388 -780 -354
rect 780 -388 876 -354
<< viali >>
rect -700 251 -492 285
rect -402 251 -194 285
rect -104 251 104 285
rect 194 251 402 285
rect 492 251 700 285
rect -762 -264 -728 192
rect -464 -264 -430 192
rect -166 -264 -132 192
rect 132 -264 166 192
rect 430 -264 464 192
rect 728 -264 762 192
<< metal1 >>
rect -712 285 -480 291
rect -712 251 -700 285
rect -492 251 -480 285
rect -712 245 -480 251
rect -414 285 -182 291
rect -414 251 -402 285
rect -194 251 -182 285
rect -414 245 -182 251
rect -116 285 116 291
rect -116 251 -104 285
rect 104 251 116 285
rect -116 245 116 251
rect 182 285 414 291
rect 182 251 194 285
rect 402 251 414 285
rect 182 245 414 251
rect 480 285 712 291
rect 480 251 492 285
rect 700 251 712 285
rect 480 245 712 251
rect -768 192 -722 204
rect -768 -264 -762 192
rect -728 -264 -722 192
rect -768 -276 -722 -264
rect -470 192 -424 204
rect -470 -264 -464 192
rect -430 -264 -424 192
rect -470 -276 -424 -264
rect -172 192 -126 204
rect -172 -264 -166 192
rect -132 -264 -126 192
rect -172 -276 -126 -264
rect 126 192 172 204
rect 126 -264 132 192
rect 166 -264 172 192
rect 126 -276 172 -264
rect 424 192 470 204
rect 424 -264 430 192
rect 464 -264 470 192
rect 424 -276 470 -264
rect 722 192 768 204
rect 722 -264 728 192
rect 762 -264 768 192
rect 722 -276 768 -264
<< properties >>
string FIXED_BBOX -859 -371 859 371
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 2.4 l 1.2 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
