magic
tech sky130A
magscale 1 2
timestamp 1663450919
<< pwell >>
rect -246 -329 246 329
<< nmoslvt >>
rect -50 -119 50 181
<< ndiff >>
rect -108 169 -50 181
rect -108 -107 -96 169
rect -62 -107 -50 169
rect -108 -119 -50 -107
rect 50 169 108 181
rect 50 -107 62 169
rect 96 -107 108 169
rect 50 -119 108 -107
<< ndiffc >>
rect -96 -107 -62 169
rect 62 -107 96 169
<< psubdiff >>
rect -210 259 -114 293
rect 114 259 210 293
rect -210 197 -176 259
rect 176 197 210 259
rect -210 -259 -176 -197
rect 176 -259 210 -197
rect -210 -293 -114 -259
rect 114 -293 210 -259
<< psubdiffcont >>
rect -114 259 114 293
rect -210 -197 -176 197
rect 176 -197 210 197
rect -114 -293 114 -259
<< poly >>
rect -50 181 50 207
rect -50 -157 50 -119
rect -50 -191 -34 -157
rect 34 -191 50 -157
rect -50 -207 50 -191
<< polycont >>
rect -34 -191 34 -157
<< locali >>
rect -210 259 -114 293
rect 114 259 210 293
rect -210 197 -176 259
rect 176 197 210 259
rect -96 169 -62 185
rect -96 -123 -62 -107
rect 62 169 96 185
rect 62 -123 96 -107
rect -50 -191 -34 -157
rect 34 -191 50 -157
rect -210 -259 -176 -197
rect 176 -259 210 -197
rect -210 -293 -114 -259
rect 114 -293 210 -259
<< viali >>
rect -96 -107 -62 169
rect 62 -107 96 169
rect -34 -191 34 -157
<< metal1 >>
rect -102 169 -56 181
rect -102 -107 -96 169
rect -62 -107 -56 169
rect -102 -119 -56 -107
rect 56 169 102 181
rect 56 -107 62 169
rect 96 -107 102 169
rect 56 -119 102 -107
rect -46 -157 46 -151
rect -46 -191 -34 -157
rect 34 -191 46 -157
rect -46 -197 46 -191
<< properties >>
string FIXED_BBOX -193 -276 193 276
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.5 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
