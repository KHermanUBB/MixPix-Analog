magic
tech sky130A
magscale 1 2
timestamp 1663448085
<< nwell >>
rect -912 -424 912 424
<< pmoslvt >>
rect -716 -204 -476 276
rect -418 -204 -178 276
rect -120 -204 120 276
rect 178 -204 418 276
rect 476 -204 716 276
<< pdiff >>
rect -774 264 -716 276
rect -774 -192 -762 264
rect -728 -192 -716 264
rect -774 -204 -716 -192
rect -476 264 -418 276
rect -476 -192 -464 264
rect -430 -192 -418 264
rect -476 -204 -418 -192
rect -178 264 -120 276
rect -178 -192 -166 264
rect -132 -192 -120 264
rect -178 -204 -120 -192
rect 120 264 178 276
rect 120 -192 132 264
rect 166 -192 178 264
rect 120 -204 178 -192
rect 418 264 476 276
rect 418 -192 430 264
rect 464 -192 476 264
rect 418 -204 476 -192
rect 716 264 774 276
rect 716 -192 728 264
rect 762 -192 774 264
rect 716 -204 774 -192
<< pdiffc >>
rect -762 -192 -728 264
rect -464 -192 -430 264
rect -166 -192 -132 264
rect 132 -192 166 264
rect 430 -192 464 264
rect 728 -192 762 264
<< nsubdiff >>
rect -876 354 -780 388
rect 780 354 876 388
rect -876 291 -842 354
rect 842 291 876 354
rect -876 -354 -842 -291
rect 842 -354 876 -291
rect -876 -388 -780 -354
rect 780 -388 876 -354
<< nsubdiffcont >>
rect -780 354 780 388
rect -876 -291 -842 291
rect 842 -291 876 291
rect -780 -388 780 -354
<< poly >>
rect -716 276 -476 302
rect -418 276 -178 302
rect -120 276 120 302
rect 178 276 418 302
rect 476 276 716 302
rect -716 -251 -476 -204
rect -716 -285 -700 -251
rect -492 -285 -476 -251
rect -716 -301 -476 -285
rect -418 -251 -178 -204
rect -418 -285 -402 -251
rect -194 -285 -178 -251
rect -418 -301 -178 -285
rect -120 -251 120 -204
rect -120 -285 -104 -251
rect 104 -285 120 -251
rect -120 -301 120 -285
rect 178 -251 418 -204
rect 178 -285 194 -251
rect 402 -285 418 -251
rect 178 -301 418 -285
rect 476 -251 716 -204
rect 476 -285 492 -251
rect 700 -285 716 -251
rect 476 -301 716 -285
<< polycont >>
rect -700 -285 -492 -251
rect -402 -285 -194 -251
rect -104 -285 104 -251
rect 194 -285 402 -251
rect 492 -285 700 -251
<< locali >>
rect -876 354 -780 388
rect 780 354 876 388
rect -876 291 -842 354
rect 842 291 876 354
rect -762 264 -728 280
rect -762 -208 -728 -192
rect -464 264 -430 280
rect -464 -208 -430 -192
rect -166 264 -132 280
rect -166 -208 -132 -192
rect 132 264 166 280
rect 132 -208 166 -192
rect 430 264 464 280
rect 430 -208 464 -192
rect 728 264 762 280
rect 728 -208 762 -192
rect -716 -285 -700 -251
rect -492 -285 -476 -251
rect -418 -285 -402 -251
rect -194 -285 -178 -251
rect -120 -285 -104 -251
rect 104 -285 120 -251
rect 178 -285 194 -251
rect 402 -285 418 -251
rect 476 -285 492 -251
rect 700 -285 716 -251
rect -876 -354 -842 -291
rect 842 -354 876 -291
rect -876 -388 -780 -354
rect 780 -388 876 -354
<< viali >>
rect -762 -192 -728 264
rect -464 -192 -430 264
rect -166 -192 -132 264
rect 132 -192 166 264
rect 430 -192 464 264
rect 728 -192 762 264
rect -700 -285 -492 -251
rect -402 -285 -194 -251
rect -104 -285 104 -251
rect 194 -285 402 -251
rect 492 -285 700 -251
<< metal1 >>
rect -768 264 -722 276
rect -768 -192 -762 264
rect -728 -192 -722 264
rect -768 -204 -722 -192
rect -470 264 -424 276
rect -470 -192 -464 264
rect -430 -192 -424 264
rect -470 -204 -424 -192
rect -172 264 -126 276
rect -172 -192 -166 264
rect -132 -192 -126 264
rect -172 -204 -126 -192
rect 126 264 172 276
rect 126 -192 132 264
rect 166 -192 172 264
rect 126 -204 172 -192
rect 424 264 470 276
rect 424 -192 430 264
rect 464 -192 470 264
rect 424 -204 470 -192
rect 722 264 768 276
rect 722 -192 728 264
rect 762 -192 768 264
rect 722 -204 768 -192
rect -712 -251 -480 -245
rect -712 -285 -700 -251
rect -492 -285 -480 -251
rect -712 -291 -480 -285
rect -414 -251 -182 -245
rect -414 -285 -402 -251
rect -194 -285 -182 -251
rect -414 -291 -182 -285
rect -116 -251 116 -245
rect -116 -285 -104 -251
rect 104 -285 116 -251
rect -116 -291 116 -285
rect 182 -251 414 -245
rect 182 -285 194 -251
rect 402 -285 414 -251
rect 182 -291 414 -285
rect 480 -251 712 -245
rect 480 -285 492 -251
rect 700 -285 712 -251
rect 480 -291 712 -285
<< properties >>
string FIXED_BBOX -859 -371 859 371
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 2.4 l 1.2 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
