magic
tech sky130A
magscale 1 2
timestamp 1663449709
<< nwell >>
rect -425 -284 425 284
<< pmoslvt >>
rect -229 -136 -29 64
rect 29 -136 229 64
<< pdiff >>
rect -287 52 -229 64
rect -287 -124 -275 52
rect -241 -124 -229 52
rect -287 -136 -229 -124
rect -29 52 29 64
rect -29 -124 -17 52
rect 17 -124 29 52
rect -29 -136 29 -124
rect 229 52 287 64
rect 229 -124 241 52
rect 275 -124 287 52
rect 229 -136 287 -124
<< pdiffc >>
rect -275 -124 -241 52
rect -17 -124 17 52
rect 241 -124 275 52
<< nsubdiff >>
rect -389 214 -293 248
rect 293 214 389 248
rect -389 151 -355 214
rect 355 151 389 214
rect -389 -214 -355 -151
rect 355 -214 389 -151
rect -389 -248 -293 -214
rect 293 -248 389 -214
<< nsubdiffcont >>
rect -293 214 293 248
rect -389 -151 -355 151
rect 355 -151 389 151
rect -293 -248 293 -214
<< poly >>
rect -229 145 -29 161
rect -229 111 -213 145
rect -45 111 -29 145
rect -229 64 -29 111
rect 29 145 229 161
rect 29 111 45 145
rect 213 111 229 145
rect 29 64 229 111
rect -229 -162 -29 -136
rect 29 -162 229 -136
<< polycont >>
rect -213 111 -45 145
rect 45 111 213 145
<< locali >>
rect -389 214 -293 248
rect 293 214 389 248
rect -389 151 -355 214
rect 355 151 389 214
rect -229 111 -213 145
rect -45 111 -29 145
rect 29 111 45 145
rect 213 111 229 145
rect -275 52 -241 68
rect -275 -140 -241 -124
rect -17 52 17 68
rect -17 -140 17 -124
rect 241 52 275 68
rect 241 -140 275 -124
rect -389 -214 -355 -151
rect 355 -214 389 -151
rect -389 -248 -293 -214
rect 293 -248 389 -214
<< viali >>
rect -213 111 -45 145
rect 45 111 213 145
rect -275 -124 -241 52
rect -17 -124 17 52
rect 241 -124 275 52
<< metal1 >>
rect -225 145 -33 151
rect -225 111 -213 145
rect -45 111 -33 145
rect -225 105 -33 111
rect 33 145 225 151
rect 33 111 45 145
rect 213 111 225 145
rect 33 105 225 111
rect -281 52 -235 64
rect -281 -124 -275 52
rect -241 -124 -235 52
rect -281 -136 -235 -124
rect -23 52 23 64
rect -23 -124 -17 52
rect 17 -124 23 52
rect -23 -136 23 -124
rect 235 52 281 64
rect 235 -124 241 52
rect 275 -124 281 52
rect 235 -136 281 -124
<< properties >>
string FIXED_BBOX -372 -231 372 231
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1 l 1 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
