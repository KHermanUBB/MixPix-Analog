magic
tech sky130A
magscale 1 2
timestamp 1663448045
<< pwell >>
rect -1457 -429 1457 429
<< nmoslvt >>
rect -1261 -281 -1061 219
rect -1003 -281 -803 219
rect -745 -281 -545 219
rect -487 -281 -287 219
rect -229 -281 -29 219
rect 29 -281 229 219
rect 287 -281 487 219
rect 545 -281 745 219
rect 803 -281 1003 219
rect 1061 -281 1261 219
<< ndiff >>
rect -1319 207 -1261 219
rect -1319 -269 -1307 207
rect -1273 -269 -1261 207
rect -1319 -281 -1261 -269
rect -1061 207 -1003 219
rect -1061 -269 -1049 207
rect -1015 -269 -1003 207
rect -1061 -281 -1003 -269
rect -803 207 -745 219
rect -803 -269 -791 207
rect -757 -269 -745 207
rect -803 -281 -745 -269
rect -545 207 -487 219
rect -545 -269 -533 207
rect -499 -269 -487 207
rect -545 -281 -487 -269
rect -287 207 -229 219
rect -287 -269 -275 207
rect -241 -269 -229 207
rect -287 -281 -229 -269
rect -29 207 29 219
rect -29 -269 -17 207
rect 17 -269 29 207
rect -29 -281 29 -269
rect 229 207 287 219
rect 229 -269 241 207
rect 275 -269 287 207
rect 229 -281 287 -269
rect 487 207 545 219
rect 487 -269 499 207
rect 533 -269 545 207
rect 487 -281 545 -269
rect 745 207 803 219
rect 745 -269 757 207
rect 791 -269 803 207
rect 745 -281 803 -269
rect 1003 207 1061 219
rect 1003 -269 1015 207
rect 1049 -269 1061 207
rect 1003 -281 1061 -269
rect 1261 207 1319 219
rect 1261 -269 1273 207
rect 1307 -269 1319 207
rect 1261 -281 1319 -269
<< ndiffc >>
rect -1307 -269 -1273 207
rect -1049 -269 -1015 207
rect -791 -269 -757 207
rect -533 -269 -499 207
rect -275 -269 -241 207
rect -17 -269 17 207
rect 241 -269 275 207
rect 499 -269 533 207
rect 757 -269 791 207
rect 1015 -269 1049 207
rect 1273 -269 1307 207
<< psubdiff >>
rect -1421 359 -1325 393
rect 1325 359 1421 393
rect -1421 297 -1387 359
rect 1387 297 1421 359
rect -1421 -359 -1387 -297
rect 1387 -359 1421 -297
rect -1421 -393 -1325 -359
rect 1325 -393 1421 -359
<< psubdiffcont >>
rect -1325 359 1325 393
rect -1421 -297 -1387 297
rect 1387 -297 1421 297
rect -1325 -393 1325 -359
<< poly >>
rect -1261 291 -1061 307
rect -1261 257 -1245 291
rect -1077 257 -1061 291
rect -1261 219 -1061 257
rect -1003 291 -803 307
rect -1003 257 -987 291
rect -819 257 -803 291
rect -1003 219 -803 257
rect -745 291 -545 307
rect -745 257 -729 291
rect -561 257 -545 291
rect -745 219 -545 257
rect -487 291 -287 307
rect -487 257 -471 291
rect -303 257 -287 291
rect -487 219 -287 257
rect -229 291 -29 307
rect -229 257 -213 291
rect -45 257 -29 291
rect -229 219 -29 257
rect 29 291 229 307
rect 29 257 45 291
rect 213 257 229 291
rect 29 219 229 257
rect 287 291 487 307
rect 287 257 303 291
rect 471 257 487 291
rect 287 219 487 257
rect 545 291 745 307
rect 545 257 561 291
rect 729 257 745 291
rect 545 219 745 257
rect 803 291 1003 307
rect 803 257 819 291
rect 987 257 1003 291
rect 803 219 1003 257
rect 1061 291 1261 307
rect 1061 257 1077 291
rect 1245 257 1261 291
rect 1061 219 1261 257
rect -1261 -307 -1061 -281
rect -1003 -307 -803 -281
rect -745 -307 -545 -281
rect -487 -307 -287 -281
rect -229 -307 -29 -281
rect 29 -307 229 -281
rect 287 -307 487 -281
rect 545 -307 745 -281
rect 803 -307 1003 -281
rect 1061 -307 1261 -281
<< polycont >>
rect -1245 257 -1077 291
rect -987 257 -819 291
rect -729 257 -561 291
rect -471 257 -303 291
rect -213 257 -45 291
rect 45 257 213 291
rect 303 257 471 291
rect 561 257 729 291
rect 819 257 987 291
rect 1077 257 1245 291
<< locali >>
rect -1421 359 -1325 393
rect 1325 359 1421 393
rect -1421 297 -1387 359
rect 1387 297 1421 359
rect -1261 257 -1245 291
rect -1077 257 -1061 291
rect -1003 257 -987 291
rect -819 257 -803 291
rect -745 257 -729 291
rect -561 257 -545 291
rect -487 257 -471 291
rect -303 257 -287 291
rect -229 257 -213 291
rect -45 257 -29 291
rect 29 257 45 291
rect 213 257 229 291
rect 287 257 303 291
rect 471 257 487 291
rect 545 257 561 291
rect 729 257 745 291
rect 803 257 819 291
rect 987 257 1003 291
rect 1061 257 1077 291
rect 1245 257 1261 291
rect -1307 207 -1273 223
rect -1307 -285 -1273 -269
rect -1049 207 -1015 223
rect -1049 -285 -1015 -269
rect -791 207 -757 223
rect -791 -285 -757 -269
rect -533 207 -499 223
rect -533 -285 -499 -269
rect -275 207 -241 223
rect -275 -285 -241 -269
rect -17 207 17 223
rect -17 -285 17 -269
rect 241 207 275 223
rect 241 -285 275 -269
rect 499 207 533 223
rect 499 -285 533 -269
rect 757 207 791 223
rect 757 -285 791 -269
rect 1015 207 1049 223
rect 1015 -285 1049 -269
rect 1273 207 1307 223
rect 1273 -285 1307 -269
rect -1421 -359 -1387 -297
rect 1387 -359 1421 -297
rect -1421 -393 -1325 -359
rect 1325 -393 1421 -359
<< viali >>
rect -1245 257 -1077 291
rect -987 257 -819 291
rect -729 257 -561 291
rect -471 257 -303 291
rect -213 257 -45 291
rect 45 257 213 291
rect 303 257 471 291
rect 561 257 729 291
rect 819 257 987 291
rect 1077 257 1245 291
rect -1307 -269 -1273 207
rect -1049 -269 -1015 207
rect -791 -269 -757 207
rect -533 -269 -499 207
rect -275 -269 -241 207
rect -17 -269 17 207
rect 241 -269 275 207
rect 499 -269 533 207
rect 757 -269 791 207
rect 1015 -269 1049 207
rect 1273 -269 1307 207
<< metal1 >>
rect -1257 291 -1065 297
rect -1257 257 -1245 291
rect -1077 257 -1065 291
rect -1257 251 -1065 257
rect -999 291 -807 297
rect -999 257 -987 291
rect -819 257 -807 291
rect -999 251 -807 257
rect -741 291 -549 297
rect -741 257 -729 291
rect -561 257 -549 291
rect -741 251 -549 257
rect -483 291 -291 297
rect -483 257 -471 291
rect -303 257 -291 291
rect -483 251 -291 257
rect -225 291 -33 297
rect -225 257 -213 291
rect -45 257 -33 291
rect -225 251 -33 257
rect 33 291 225 297
rect 33 257 45 291
rect 213 257 225 291
rect 33 251 225 257
rect 291 291 483 297
rect 291 257 303 291
rect 471 257 483 291
rect 291 251 483 257
rect 549 291 741 297
rect 549 257 561 291
rect 729 257 741 291
rect 549 251 741 257
rect 807 291 999 297
rect 807 257 819 291
rect 987 257 999 291
rect 807 251 999 257
rect 1065 291 1257 297
rect 1065 257 1077 291
rect 1245 257 1257 291
rect 1065 251 1257 257
rect -1313 207 -1267 219
rect -1313 -269 -1307 207
rect -1273 -269 -1267 207
rect -1313 -281 -1267 -269
rect -1055 207 -1009 219
rect -1055 -269 -1049 207
rect -1015 -269 -1009 207
rect -1055 -281 -1009 -269
rect -797 207 -751 219
rect -797 -269 -791 207
rect -757 -269 -751 207
rect -797 -281 -751 -269
rect -539 207 -493 219
rect -539 -269 -533 207
rect -499 -269 -493 207
rect -539 -281 -493 -269
rect -281 207 -235 219
rect -281 -269 -275 207
rect -241 -269 -235 207
rect -281 -281 -235 -269
rect -23 207 23 219
rect -23 -269 -17 207
rect 17 -269 23 207
rect -23 -281 23 -269
rect 235 207 281 219
rect 235 -269 241 207
rect 275 -269 281 207
rect 235 -281 281 -269
rect 493 207 539 219
rect 493 -269 499 207
rect 533 -269 539 207
rect 493 -281 539 -269
rect 751 207 797 219
rect 751 -269 757 207
rect 791 -269 797 207
rect 751 -281 797 -269
rect 1009 207 1055 219
rect 1009 -269 1015 207
rect 1049 -269 1055 207
rect 1009 -281 1055 -269
rect 1267 207 1313 219
rect 1267 -269 1273 207
rect 1307 -269 1313 207
rect 1267 -281 1313 -269
<< properties >>
string FIXED_BBOX -1404 -376 1404 376
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2.5 l 1.0 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
