magic
tech sky130A
magscale 1 2
timestamp 1663448021
<< nwell >>
rect -296 -731 296 731
<< pmoslvt >>
rect -100 -512 100 512
<< pdiff >>
rect -158 500 -100 512
rect -158 -500 -146 500
rect -112 -500 -100 500
rect -158 -512 -100 -500
rect 100 500 158 512
rect 100 -500 112 500
rect 146 -500 158 500
rect 100 -512 158 -500
<< pdiffc >>
rect -146 -500 -112 500
rect 112 -500 146 500
<< nsubdiff >>
rect -260 661 -164 695
rect 164 661 260 695
rect -260 599 -226 661
rect 226 599 260 661
rect -260 -661 -226 -599
rect 226 -661 260 -599
rect -260 -695 -164 -661
rect 164 -695 260 -661
<< nsubdiffcont >>
rect -164 661 164 695
rect -260 -599 -226 599
rect 226 -599 260 599
rect -164 -695 164 -661
<< poly >>
rect -100 593 100 609
rect -100 559 -84 593
rect 84 559 100 593
rect -100 512 100 559
rect -100 -559 100 -512
rect -100 -593 -84 -559
rect 84 -593 100 -559
rect -100 -609 100 -593
<< polycont >>
rect -84 559 84 593
rect -84 -593 84 -559
<< locali >>
rect -260 661 -164 695
rect 164 661 260 695
rect -260 599 -226 661
rect 226 599 260 661
rect -100 559 -84 593
rect 84 559 100 593
rect -146 500 -112 516
rect -146 -516 -112 -500
rect 112 500 146 516
rect 112 -516 146 -500
rect -100 -593 -84 -559
rect 84 -593 100 -559
rect -260 -661 -226 -599
rect 226 -661 260 -599
rect -260 -695 -164 -661
rect 164 -695 260 -661
<< viali >>
rect -84 559 84 593
rect -146 -500 -112 500
rect 112 -500 146 500
rect -84 -593 84 -559
<< metal1 >>
rect -96 593 96 599
rect -96 559 -84 593
rect 84 559 96 593
rect -96 553 96 559
rect -152 500 -106 512
rect -152 -500 -146 500
rect -112 -500 -106 500
rect -152 -512 -106 -500
rect 106 500 152 512
rect 106 -500 112 500
rect 146 -500 152 500
rect 106 -512 152 -500
rect -96 -559 96 -553
rect -96 -593 -84 -559
rect 84 -593 96 -559
rect -96 -599 96 -593
<< properties >>
string FIXED_BBOX -243 -678 243 678
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 5.12 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
