magic
tech sky130A
timestamp 1663448021
<< pwell >>
rect -148 -1355 148 1355
<< nmoslvt >>
rect -50 -1250 50 1250
<< ndiff >>
rect -79 1244 -50 1250
rect -79 -1244 -73 1244
rect -56 -1244 -50 1244
rect -79 -1250 -50 -1244
rect 50 1244 79 1250
rect 50 -1244 56 1244
rect 73 -1244 79 1244
rect 50 -1250 79 -1244
<< ndiffc >>
rect -73 -1244 -56 1244
rect 56 -1244 73 1244
<< psubdiff >>
rect -130 1320 -82 1337
rect 82 1320 130 1337
rect -130 1289 -113 1320
rect 113 1289 130 1320
rect -130 -1320 -113 -1289
rect 113 -1320 130 -1289
rect -130 -1337 -82 -1320
rect 82 -1337 130 -1320
<< psubdiffcont >>
rect -82 1320 82 1337
rect -130 -1289 -113 1289
rect 113 -1289 130 1289
rect -82 -1337 82 -1320
<< poly >>
rect -50 1286 50 1294
rect -50 1269 -42 1286
rect 42 1269 50 1286
rect -50 1250 50 1269
rect -50 -1269 50 -1250
rect -50 -1286 -42 -1269
rect 42 -1286 50 -1269
rect -50 -1294 50 -1286
<< polycont >>
rect -42 1269 42 1286
rect -42 -1286 42 -1269
<< locali >>
rect -130 1320 -82 1337
rect 82 1320 130 1337
rect -130 1289 -113 1320
rect 113 1289 130 1320
rect -50 1269 -42 1286
rect 42 1269 50 1286
rect -73 1244 -56 1252
rect -73 -1252 -56 -1244
rect 56 1244 73 1252
rect 56 -1252 73 -1244
rect -50 -1286 -42 -1269
rect 42 -1286 50 -1269
rect -130 -1320 -113 -1289
rect 113 -1320 130 -1289
rect -130 -1337 -82 -1320
rect 82 -1337 130 -1320
<< viali >>
rect -42 1269 42 1286
rect -73 -1244 -56 1244
rect 56 -1244 73 1244
rect -42 -1286 42 -1269
<< metal1 >>
rect -48 1286 48 1289
rect -48 1269 -42 1286
rect 42 1269 48 1286
rect -48 1266 48 1269
rect -76 1244 -53 1250
rect -76 -1244 -73 1244
rect -56 -1244 -53 1244
rect -76 -1250 -53 -1244
rect 53 1244 76 1250
rect 53 -1244 56 1244
rect 73 -1244 76 1244
rect 53 -1250 76 -1244
rect -48 -1269 48 -1266
rect -48 -1286 -42 -1269
rect 42 -1286 48 -1269
rect -48 -1289 48 -1286
<< properties >>
string FIXED_BBOX -121 -1328 121 1328
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 25.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
