** sch_path: /home/krzysztof/asic/analog/nmos_characterization/nmos3_3.sch
**.subckt nmos3_3
VDD net1 GND 1.8
Vg net2 GND 0
Vm net3 net1 0
XM1 net3 net2 GND GND sky130_fd_pr__nfet_01v8_lvt L={L} W={W} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code
** opencircuitdesign pdks install
.lib /home/icarosix/asic/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
**** end user architecture code
**.ends
.GLOBAL GND
**** begin user architecture code
* .option SCALE=1e-6
.option method=gear seed=12
.param L=2
.param W=1
.DC Vg 0.2 0.7 0.001
.control
set hcopydevtype = svg
set nolegend
set color0=white
set color1=black
set color2=blue
set color3=red
*****************************************************************************
 run
let Vgs = V(net2)
let Id = -vm#branch
let gm_id = deriv(Id)/Id 
save all
write all
meas dc Vgs2 when gm_id=10
meas dc  Id2 find Id when  Vgs=Vgs2
*hardcopy IDoutput.svg xlabel "Vds" ylabel "Id" title "Drian current"  -I(Vm)
 plot xlabel "Vgs" ylabel "gm/Id" title "Gm over ID"   deriv(Id)/Id 
* plot   -I(Vm)
*hardcopy gm_ID.svg xlabel "Vgs" ylabel "Id" title "Drian current"  -I(Vm)
*hardcopy gmoverID_vsVgs.svg    xlabel "Vgs" ylabel "gm/Id" title "Gm over ID"   deriv(I(Vm))/I(Vm)
******************************************************************************
.endc
.end
