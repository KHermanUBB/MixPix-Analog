../xchem/simulation/OTA3_kh_PVersion.spice