magic
tech sky130A
magscale 1 2
timestamp 1663448021
<< nwell >>
rect -316 -1419 316 1419
<< pmoslvt >>
rect -120 -1200 120 1200
<< pdiff >>
rect -178 1188 -120 1200
rect -178 -1188 -166 1188
rect -132 -1188 -120 1188
rect -178 -1200 -120 -1188
rect 120 1188 178 1200
rect 120 -1188 132 1188
rect 166 -1188 178 1188
rect 120 -1200 178 -1188
<< pdiffc >>
rect -166 -1188 -132 1188
rect 132 -1188 166 1188
<< nsubdiff >>
rect -280 1349 -184 1383
rect 184 1349 280 1383
rect -280 1287 -246 1349
rect 246 1287 280 1349
rect -280 -1349 -246 -1287
rect 246 -1349 280 -1287
rect -280 -1383 -184 -1349
rect 184 -1383 280 -1349
<< nsubdiffcont >>
rect -184 1349 184 1383
rect -280 -1287 -246 1287
rect 246 -1287 280 1287
rect -184 -1383 184 -1349
<< poly >>
rect -120 1281 120 1297
rect -120 1247 -104 1281
rect 104 1247 120 1281
rect -120 1200 120 1247
rect -120 -1247 120 -1200
rect -120 -1281 -104 -1247
rect 104 -1281 120 -1247
rect -120 -1297 120 -1281
<< polycont >>
rect -104 1247 104 1281
rect -104 -1281 104 -1247
<< locali >>
rect -280 1349 -184 1383
rect 184 1349 280 1383
rect -280 1287 -246 1349
rect 246 1287 280 1349
rect -120 1247 -104 1281
rect 104 1247 120 1281
rect -166 1188 -132 1204
rect -166 -1204 -132 -1188
rect 132 1188 166 1204
rect 132 -1204 166 -1188
rect -120 -1281 -104 -1247
rect 104 -1281 120 -1247
rect -280 -1349 -246 -1287
rect 246 -1349 280 -1287
rect -280 -1383 -184 -1349
rect 184 -1383 280 -1349
<< viali >>
rect -104 1247 104 1281
rect -166 -1188 -132 1188
rect 132 -1188 166 1188
rect -104 -1281 104 -1247
<< metal1 >>
rect -116 1281 116 1287
rect -116 1247 -104 1281
rect 104 1247 116 1281
rect -116 1241 116 1247
rect -172 1188 -126 1200
rect -172 -1188 -166 1188
rect -132 -1188 -126 1188
rect -172 -1200 -126 -1188
rect 126 1188 172 1200
rect 126 -1188 132 1188
rect 166 -1188 172 1188
rect 126 -1200 172 -1188
rect -116 -1247 116 -1241
rect -116 -1281 -104 -1247
rect 104 -1281 116 -1247
rect -116 -1287 116 -1281
<< properties >>
string FIXED_BBOX -263 -1366 263 1366
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 12.0 l 1.2 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
